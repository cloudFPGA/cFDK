module Hash
(
    Key,
    Hash
);

// lookup parameters
localparam K = 97; // number of key bits
localparam H = 48; // number of hash bits

// I/O declarations
input   [K-1:0]     Key;
output  [H-1:0]     Hash;

//*************************************
reg     [H-1:0]     Hash;

// calculate hash
always @* begin
    Hash[0] = ^{ Key & 97'b1011010111000011111110111000110000010111001100110111010000100001111001101110101110101100101110100 };
    Hash[1] = ^{ Key & 97'b0011001110111000111110100100101001111110101110000010010101010110010011000010001000110101101110010 };
    Hash[2] = ^{ Key & 97'b1101100111100111111010101100110101010001110100010001101011110111110111110110010011100011110000000 };
    Hash[3] = ^{ Key & 97'b0100111010110001111000010101000010101100111000000000110010000000100001111100101111101110110111100 };
    Hash[4] = ^{ Key & 97'b0100101001000101100111100110100110111101010001101011110000001000011001100110011011111100110101111 };
    Hash[5] = ^{ Key & 97'b0011100111010101000001100011010000010101110000110010001100001010101000011101001101010110101001010 };
    Hash[6] = ^{ Key & 97'b1000001100010100000001001100111111010011010011101100100011111111101000110101001100110011011101011 };
    Hash[7] = ^{ Key & 97'b1011001111100010111010001110010111010111100111001000100011011011000101011100001011110110011001111 };
    Hash[8] = ^{ Key & 97'b0110110101001111110011110100000111111010011000011101001100111111100000001011000100110110101010101 };
    Hash[9] = ^{ Key & 97'b1101001100011101101100001011100011001110011111001101000001011000101010011001100000110001001111110 };
    Hash[10] = ^{ Key & 97'b0011110100101010000000011111110001011010011100001011110100010101001011100001000001111000001100110 };
    Hash[11] = ^{ Key & 97'b0110111100101000000011110111110110010010110010001101111010001101001110011001110110000000000001010 };
    Hash[12] = ^{ Key & 97'b0011001001011101101100111001111000100100101101100001101111111010001100001001110110000001001001111 };
    Hash[13] = ^{ Key & 97'b1010011111011101100010101110011000001010100010111100110001010111110010110011000001001010000000110 };
    Hash[14] = ^{ Key & 97'b0010010101100000110110100110001111110101001101101011001101100100001011100111010101001000011100011 };
    Hash[15] = ^{ Key & 97'b1101110011000011011000111010011011111110011100000000000011101111111100101011111100100001010100101 };
    Hash[16] = ^{ Key & 97'b0110001011010110000100001111001110111111011101010111110100011000101100000010111011000110000111000 };
    Hash[17] = ^{ Key & 97'b1110010101111010100110011101011100000100101010001111010010101110010011110100010110010101001011110 };
    Hash[18] = ^{ Key & 97'b0011011111101010110110000011110110001001000010100001011111111110001110111000110010001110111100111 };
    Hash[19] = ^{ Key & 97'b1000100100110000110101000010011001100000001011111011101000010001011001000110001111101001101111001 };
    Hash[20] = ^{ Key & 97'b1001001100110001000000101101111011001100100000010110110011000001010011000000001100001101110010100 };
    Hash[21] = ^{ Key & 97'b1101001011011110101011001001001010111010010100000100110111000010011101110110101010010000111101101 };
    Hash[22] = ^{ Key & 97'b1110101010101000111011110100001000100011010011110110001110011001000001000010110011001001111111010 };
    Hash[23] = ^{ Key & 97'b1110000011111100010011101111100100001111010111100000101101010101110001010001100001111101111100100 };
    Hash[24] = ^{ Key & 97'b0001001001000101010010011001111111100011110010101101110010100000111110110010001001110011100111001 };
    Hash[25] = ^{ Key & 97'b0111111010101010001101000011111101000011100101110011000110101010011011111101010111011000011111100 };
    Hash[26] = ^{ Key & 97'b0000100010010010010001001101001100110011101100010010010100001010000111001001111110111110101010011 };
    Hash[27] = ^{ Key & 97'b0010111000110010000111010101100100011110110010011100110111101000101001101100110001110011100100001 };
    Hash[28] = ^{ Key & 97'b0111001010100001101011101011000101000101001111101100000011100101010010101111100100010110110111101 };
    Hash[29] = ^{ Key & 97'b1100110110000111000100011010001011000101111101100111001100111000010100000100100110111010001111011 };
    Hash[30] = ^{ Key & 97'b1000110000001110111111111001010001001000001001101110001000111101000101010111011001100011010000010 };
    Hash[31] = ^{ Key & 97'b1110010001001001000001110010010111100001100100001100111001100011110111001011011000000001011011001 };
    Hash[32] = ^{ Key & 97'b1001111001011101011101111011111111011111000110110011011001111010001000101000111001110101100010001 };
    Hash[33] = ^{ Key & 97'b0000001100111011001101010111100000101000101000111001001010111100101110011111110010011101100010100 };
    Hash[34] = ^{ Key & 97'b1101010100110111001111011000110110110000110100110011111110001101110000010111111100111100010001001 };
    Hash[35] = ^{ Key & 97'b1001110101001100001101010110110111011010000011011111111101001100000010010100001110001001110110010 };
    Hash[36] = ^{ Key & 97'b1110010101000100110001010001101101011001100111000010001100000111000101001100110001011111001000110 };
    Hash[37] = ^{ Key & 97'b0100000110010100011010111011001100011101111110011010000111101110010111111011000111000010010111111 };
    Hash[38] = ^{ Key & 97'b1110101010101000011100100010010010110111011011011101110101010111110110100011001011000100110001010 };
    Hash[39] = ^{ Key & 97'b0100011000100111111101000000100000101101101111010110101010111101110111000001111100001110010011001 };
    Hash[40] = ^{ Key & 97'b0111000111010000010110110000010000100000000111110011100100100000001100000110100011000010000000100 };
    Hash[41] = ^{ Key & 97'b0001100001001011101101010101101000100001110001111100000011110001111111001101100011101101111001101 };
    Hash[42] = ^{ Key & 97'b1011011000101010010010101011011011001110010011000000101100000110011110000010000000011011000010110 };
    Hash[43] = ^{ Key & 97'b0001100011110101001110110000100011110101011001000011011010010011100110111101011101101010000010000 };
    Hash[44] = ^{ Key & 97'b1000100010011111101100100110101001101000101101100110010000110000110000111100111111000111110110001 };
    Hash[45] = ^{ Key & 97'b0111110010100111111000000100001100100010011001111100101111000111100110111010011110001101001000011 };
    Hash[46] = ^{ Key & 97'b1000111110111110100001011000000010001000100010011100011111010011101000111001100100111110010101001 };
    Hash[47] = ^{ Key & 97'b0101110001011011010011000100001111110110001010111001011001100110111101110010010000110011101000110 };
end

//*************************************

endmodule
