fab@bivio.zurich.ibm.com.11750:1619949767