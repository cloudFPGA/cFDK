// *****************************************************************************
// *
// *                             cloudFPGA
// *            All rights reserved -- Property of IBM
// *
// *----------------------------------------------------------------------------
// *
// * Title : Flash version of the the 10G Ethernet I/F instantiated by the SHELL. 
// *
// * File    : tenGigEth_Flash.v
// *
// * Created : Dec. 2017
// * Authors : Francois Abel <fab@zurich.ibm.com>
// *
// * Devices : xcku060-ffva1156-2-i
// * Tools   : Vivado v2016.4 (64-bit)
// * Depends : None
// *
// * Description : This is the toplevel design for the 10 Gigabit Ethernet I/F
// *    instantiated by the shell of the FMKU2595 module equipped with a XCKU60
// *    device. It is referred to as the Flash version because it integrates a  
// *    loopback turn between the network layers L2 and L3 of the ETH0 interface.
// *    When this loopback is enabled, the data output by the AXI4-S interface
// *    of ETH0 are passed back to the AXI4-S input of the same ETH0. Otherwise,
// *    this module is neutral and data pass through it untouched.  
// * 
// * Parameters:
// *
// * Comments:
// *
// *****************************************************************************


// *****************************************************************************
// **  MODULE - 10G ETHERNET WITH LOOPBACK TURN
// *****************************************************************************

module TenGigEth_Flash (

  //-- Clocks and Resets inputs ------------------
  input             piTOP_156_25Clk,    // Freerunning
  input             piCLKT_Gt_RefClk_n,
  input             piCLKT_Gt_RefClk_p,
  input             piTOP_Reset,

  //-- Clocks and Resets outputs -----------------
  output            poETH0_CoreClk,

  //-- MMIO : Ctrl inputs and Status outputs -----
  input             piMMIO_Eth0_RxEqualizerMode,
  input             piMMIO_Eth0_PcsLoopbackEn,
  input             piMMIO_Eth0_MacLoopbackEn,
  output            poETH0_Mmio_CoreReady,
  output            poETH0_Mmio_QpllLock,
  output            poETH0_Mmio_ResetDone,    // [FIXME w/ wee]

  //-- ECON : Gigabit Transceivers ---------------
  input             piECON_Eth0_Gt_n,
  input             piECON_Eth0_Gt_p,
  output            poETH0_Econ_Gt_n,
  output            poETH0_Econ_Gt_p,
   
  //-- AXI4 Tx Stream Interface ------------------
  input     [63:0]  piLY3_Axis_tdata,
  input     [7:0]   piLY3_Axis_tkeep,
  input             piLY3_Axis_tvalid,
  input             piLY3_Axis_tlast,
  output            poLy3_Axis_tready,
  
  //-- AXI4 Rx Stream Interface ------------------  
  output     [63:0] poLy3_Axis_tdata,
  output     [7:0]  poLy3_Axis_tkeep,
  output            poLy3_Axis_tvalid,
  output            poLy3_Axis_tlast,
  input             piLY3_Axis_tready
  
  ); // End of PortList
   
// *****************************************************************************


  //============================================================================
  //  SIGNAL DECLARATIONS
  //============================================================================

  //-- Clocks ------------------------------------
  wire        sETH0_CoreClk;  // Generated by the ETH core. 
                              // Use it to clock the TX datapath.

  //-- AXI4 Stream ETH0 < -> NTS0 -----------------
  wire [63:0] sETH0_Elp_Axis_tdata,  sELP0_Eth_Axis_tdata;
  wire [ 7:0] sETH0_Elp_Axis_tkeep,  sELP0_Eth_Axis_tkeep;
  wire        sETH0_Elp_Axis_tvalid, sELP0_Eth_Axis_tvalid;
  wire        sETH0_Elp_Axis_tlast,  sELP0_Eth_Axis_tlast;
  wire        sELP0_Eth_Axis_tready, sETH0_Elp_Axis_tready;
    
  //-- End of signal declarations ---------------


  //============================================================================
  //  INST: 10G ETHERNET SUBSYSTEM (OSI Network Layers 1+2)
  //============================================================================
  TenGigEth ETH0 (
    
    //-- Clocks and Resets inputs ----------------
    .piTOP_156_25Clk              (piTOP_156_25Clk),    // Freerunning
    .piCLKT_Gt_RefClk_n           (piCLKT_Gt_RefClk_n),
    .piCLKT_Gt_RefClk_p           (piCLKT_Gt_RefClk_p),
    .piTOP_Reset                  (piTOP_Reset),
      
    //-- Clocks and Resets outputs ---------------
    .poETH0_CoreClk               (sETH0_CoreClk),
       
    //-- MMIO : Control inputs and Status outputs 
    .piMMIO_Eth0_RxEqualizerMode  (piMMIO_Eth0_RxEqualizerMode),
    .piMMIO_Eth0_PcsLoopbackEn    (piMMIO_Eth0_PcsLoopbackEn),
    .piMMIO_Eth0_MacLoopbackEn    (piMMIO_Eth0_MacLoopbackEn),
    .poETH0_Mmio_CoreReady        (poETH0_Mmio_CoreReady),
    .poETH0_Mmio_QpllLock         (poETH0_Mmio_QpllLock),
    .poETH0_Mmio_ResetDone        (/* network_init */), // [FIXME]

    //-- ECON : Gigabit Transceivers -------------
    .piECON_Eth0_Gt_n             (piECON_Eth0_Gt_n),
    .piECON_Eth0_Gt_p             (piECON_Eth0_Gt_p),
    .poETH0_Econ_Gt_n             (poETH0_Econ_Gt_n),
    .poETH0_Econ_Gt_p             (poETH0_Econ_Gt_p),
         
    //-- AXI4 Input Stream Interface -------------
    .piLY3_Axis_tdata             (sELP0_Eth_Axis_tdata),
    .piLY3_Axis_tkeep             (sELP0_Eth_Axis_tkeep),
    .piLY3_Axis_tvalid            (sELP0_Eth_Axis_tvalid),
    .piLY3_Axis_tlast             (sELP0_Eth_Axis_tlast),
    .poLy3_Axis_tready            (sETH0_Elp_Axis_tready),

    //-- AXI4 Output Stream Interface ------------  
    .poLy3_Axis_tdata             (sETH0_Elp_Axis_tdata),
    .poLy3_Axis_tkeep             (sETH0_Elp_Axis_tkeep),
    .poLy3_Axis_tvalid            (sETH0_Elp_Axis_tvalid),
    .poLy3_Axis_tlast             (sETH0_Elp_Axis_tlast),
    .piLY3_Axis_tready            (sELP0_Eth_Axis_tready)
    
  );
    

  //============================================================================
  //  INST: ETHERNET LOOPBACK TURN
  //============================================================================
  TenGigEth_Loop ELP0 (
      
        //-- Clocks and Resets inputs ------------
        .piEthCoreClk           (sETH0_CoreClk),
        .piReset_a              (piTOP_Reset),
      
        // -- MMIO : Ctrl Inp and Status Out -----
        .piLoopbackEn           (piMMIO_Eth0_MacLoopbackEn),

        //-- AXI4 Input Stream from L2 -----------
        .piLY2_Axis_tdata       (sETH0_Elp_Axis_tdata),
        .piLY2_Axis_tkeep       (sETH0_Elp_Axis_tkeep),
        .piLY2_Axis_tlast       (sETH0_Elp_Axis_tlast),
        .piLY2_Axis_tvalid      (sETH0_Elp_Axis_tvalid),
        .poLy2_Axis_tready      (sELP0_Eth_Axis_tready),
        
        //-- AXI4 Output Stream to L2 ------------
        .piLY2_Axis_tready      (sETH0_Elp_Axis_tready),
        .poLy2_Axis_tdata       (sELP0_Eth_Axis_tdata),
        .poLy2_Axis_tkeep       (sELP0_Eth_Axis_tkeep),
        .poLy2_Axis_tlast       (sELP0_Eth_Axis_tlast),
        .poLy2_Axis_tvalid      (sELP0_Eth_Axis_tvalid),
        
        //-- AXI4 Input Stream from L3 -----------
        .piLY3_Axis_tdata       (piLY3_Axis_tdata),
        .piLY3_Axis_tkeep       (piLY3_Axis_tkeep),
        .piLY3_Axis_tlast       (piLY3_Axis_tlast),
        .piLY3_Axis_tvalid      (piLY3_Axis_tvalid),        
        .poLy3_Axis_tready      (poLy3_Axis_tready),
        
        //-- AXI4 Output Stream to L3 ------------
        .piLY3_Axis_tready      (piLY3_Axis_tready),
        .poLy3_Axis_tdata       (poLy3_Axis_tdata),
        .poLy3_Axis_tkeep       (poLy3_Axis_tkeep),
        .poLy3_Axis_tlast       (poLy3_Axis_tlast),
        .poLy3_Axis_tvalid      (poLy3_Axis_tvalid)
                      
      );


  //============================================================================
  //  COMB: CONTINUOUS OUTPUT PORT ASSIGNMENTS
  //============================================================================
  assign poETH0_CoreClk = sETH0_CoreClk;

endmodule
