//                              -*- Mode: Verilog -*-
// *****************************************************************************
// *
// *                             cloudFPGA
// *            All rights reserved -- Property of IBM
// *
// *----------------------------------------------------------------------------
// *
// * Title : TCP Application Register Slice (TARS)
// *
// * Created : Apr. 2020
// * Authors : Francois Abel <fab@zurich.ibm.com>
// *
// * Tools   : Vivado v2016.4 (64-bit)
// * Depends : None
// *
// * Description : A placeholder containing the Axis Register Slice (ARS) 
// *    components involved in the TCP application interface of the Network
// *    Transport Stack (NTS). The use of such an Axis register slice is not
// *    a prerequisit but it is used here to provide timing isolation and to
// *    ease the place and routing phase.
// *
// *          +-----+     +----+     +---+
// *          |     <-----+    <-----+   |
// *          | NTS |     |TARS|     |APP|
// *          |     +----->    +----->   |
// *          +-----+     +----+     +---+
// *
// *****************************************************************************

`timescale 1ns / 1ps

// *****************************************************************************
// **  MODULE - TCP APPLICATION REGISTER SLICE
// *****************************************************************************

module TcpApplicationRegisterSlice

(

  //------------------------------------------------------
  //-- This is typically the Global Clock used all over the SHELL
  //------------------------------------------------------ 
  input          piClk,
  
  //------------------------------------------------------
  //-- This is typically the Global Reset used by the entire SHELL
  //--  or the OSI-Layer-5 reset generated by the MMIO. 
  //------------------------------------------------------ 
  input          piRst,
   
  //------------------------------------------------------
  //-- APP / Tcp / Tx Data Interfaces (.i.e TARS<-->APP)
  //------------------------------------------------------
  //---- Axis4-Stream TCP Data ---------------
  input  [ 63:0]  siAPP_Tcp_Data_tdata,
  input  [  7:0]  siAPP_Tcp_Data_tkeep,
  input           siAPP_Tcp_Data_tlast,
  input           siAPP_Tcp_Data_tvalid,
  output          siAPP_Tcp_Data_tready,
  //---- Axis4-Stream TCP Metadata -----------
  input  [ 15:0]  siAPP_Tcp_Meta_tdata,
  input           siAPP_Tcp_Meta_tvalid,
  output          siAPP_Tcp_Meta_tready,
 //---- Axis4-Stream TCP Data Status --------
  output [ 23:0]  soAPP_Tcp_DSts_tdata,
  output          soAPP_Tcp_DSts_tvalid,
  input           soAPP_Tcp_DSts_tready,
  
  //------------------------------------------------------
  //-- APP / Tcp / Rx Data Interfaces (.i.e TARS<-->APP)
  //------------------------------------------------------
  //-- Axis4-Stream TCP Data -----------------
  output [ 63:0]  soAPP_Tcp_Data_tdata,
  output [  7:0]  soAPP_Tcp_Data_tkeep,
  output          soAPP_Tcp_Data_tlast,
  output          soAPP_Tcp_Data_tvalid,
  input           soAPP_Tcp_Data_tready,
  //--  Axis4-Stream TCP Metadata ------------
  output [ 15:0]  soAPP_Tcp_Meta_tdata,
  output          soAPP_Tcp_Meta_tvalid,
  input           soAPP_Tcp_Meta_tready,
  //--  Axis4-Stream TCP Data Notification ---
  output [103:0]  soAPP_Tcp_Notif_tdata,  // 7+96
  output          soAPP_Tcp_Notif_tvalid,
  input           soAPP_Tcp_Notif_tready,
   //--  Axis4-Stream TCP Data Request --------
  input  [ 31:0]  siAPP_Tcp_DReq_tdata,
  input           siAPP_Tcp_DReq_tvalid,
  output          siAPP_Tcp_DReq_tready,

  //------------------------------------------------------
  //-- APP / Tcp / Tx Ctlr Interfaces (.i.e TARS<-->APP)
  //------------------------------------------------------
  //---- Axis4-Stream TCP Open Session Request
  input [ 47:0]  siAPP_Tcp_OpnReq_tdata,
  input          siAPP_Tcp_OpnReq_tvalid,
  output         siAPP_Tcp_OpnReq_tready,
  //---- Axis4-Stream TCP Open Session Reply
  output [ 23:0] soAPP_Tcp_OpnRep_tdata,
  output         soAPP_Tcp_OpnRep_tvalid,
  input          soAPP_Tcp_OpnRep_tready,
  //---- Axis4-Stream TCP Close Request ------
  input [ 15:0]  siAPP_Tcp_ClsReq_tdata,
  input          siAPP_Tcp_ClsReq_tvalid,
  output         siAPP_Tcp_ClsReq_tready,

  //------------------------------------------------------
  //-- APP / Tcp / Rx Ctlr Interfaces (.i.e TARS<-->APP)
  //------------------------------------------------------
  //----  Axis4-Stream TCP Listen Request ----
  input [ 15:0]  siAPP_Tcp_LsnReq_tdata,   
  input          siAPP_Tcp_LsnReq_tvalid,
  output         siAPP_Tcp_LsnReq_tready,
  //----  Axis4-Stream TCP Listen Rep --------
  output [  7:0] soAPP_Tcp_LsnRep_tdata,
  output         soAPP_Tcp_LsnRep_tvalid,
  input          soAPP_Tcp_LsnRep_tready,
  
  //------------------------------------------------------
  //-- NTS / Tcp / Tx Data Interfaces (.i.e NTS<-->TARS)
  //------------------------------------------------------
  //---- Axis4-Stream TCP Data ---------------
  output [ 63:0]  soNTS_Tcp_Data_tdata,
  output [  7:0]  soNTS_Tcp_Data_tkeep,
  output          soNTS_Tcp_Data_tlast,
  output          soNTS_Tcp_Data_tvalid,
  input           soNTS_Tcp_Data_tready,
  //---- Axis4-Stream TCP Metadata -----------
  output [ 15:0]  soNTS_Tcp_Meta_tdata,
  output          soNTS_Tcp_Meta_tvalid,
  input           soNTS_Tcp_Meta_tready,
  //---- Axis4-Stream TCP Data Status --------
  input  [ 23:0]  siNTS_Tcp_DSts_tdata,
  input           siNTS_Tcp_DSts_tvalid,
  output          siNTS_Tcp_DSts_tready,
    
  //------------------------------------------------------
  //-- NTS / Tcp / Rx Data Interfaces (.i.e NTS<-->TARS)
  //------------------------------------------------------
  //-- Axis4-Stream TCP Data -----------------
  input  [ 63:0]  siNTS_Tcp_Data_tdata,
  input  [  7:0]  siNTS_Tcp_Data_tkeep,
  input           siNTS_Tcp_Data_tlast,
  input           siNTS_Tcp_Data_tvalid,
  output          siNTS_Tcp_Data_tready,
  //--  Axis4-Stream TCP Metadata ------------
  input  [ 15:0]  siNTS_Tcp_Meta_tdata,
  input           siNTS_Tcp_Meta_tvalid,
  output          siNTS_Tcp_Meta_tready,
  //--  Axis4-Stream TCP Data Notification ---
  input  [103:0]  siNTS_Tcp_Notif_tdata,  // 7+96
  input           siNTS_Tcp_Notif_tvalid,
  output          siNTS_Tcp_Notif_tready,
  //--  Axis4-Stream TCP Data Request --------
  output [ 31:0]  soNTS_Tcp_DReq_tdata,
  output          soNTS_Tcp_DReq_tvalid,
  input           soNTS_Tcp_DReq_tready,
  
  //------------------------------------------------------
  //-- NTS / Tcp / Tx Ctlr Interfaces (.i.e NTS<-->TARS)
  //------------------------------------------------------
  //---- Axis4-Stream TCP Open Session Request
  output[ 47:0]  soNTS_Tcp_OpnReq_tdata,
  output         soNTS_Tcp_OpnReq_tvalid,
  input          soNTS_Tcp_OpnReq_tready,
  //---- Axis4-Stream TCP Open Session Reply
  input  [ 23:0] siNTS_Tcp_OpnRep_tdata,
  input          siNTS_Tcp_OpnRep_tvalid,
  output         siNTS_Tcp_OpnRep_tready,
  //---- Axis4-Stream TCP Close Request ------
  output[ 15:0]  soNTS_Tcp_ClsReq_tdata,
  output         soNTS_Tcp_ClsReq_tvalid,
  input          soNTS_Tcp_ClsReq_tready,
  
  //------------------------------------------------------
  //-- NTS / Tcp / Rx Ctlr Interfaces (.i.e NTS<-->TARS)
  //------------------------------------------------------
  //----  Axis4-Stream TCP Listen Request ----
  output[ 15:0]  soNTS_Tcp_LsnReq_tdata,   
  output         soNTS_Tcp_LsnReq_tvalid,
  input          soNTS_Tcp_LsnReq_tready,
  //----  Axis4-Stream TCP Listen Rep --------
  input  [  7:0] siNTS_Tcp_LsnRep_tdata,
  input          siNTS_Tcp_LsnRep_tvalid,
  output         siNTS_Tcp_LsnRep_tready

);  // End of PortList


  // *****************************************************************************
  // **  STRUCTURE
  // *****************************************************************************

  //------------------------------------------------------
  //-- TAIF / Tx Data Interfaces
  //------------------------------------------------------
  AxisRegisterSlice_64 APP_NTS_Tcp_Data (
    .aclk           (piClk),
    .aresetn        (~piRst),
    //-- From APP ----------------------
    .s_axis_tdata   (siAPP_Tcp_Data_tdata),
    .s_axis_tvalid  (siAPP_Tcp_Data_tvalid),
    .s_axis_tkeep   (siAPP_Tcp_Data_tkeep),
    .s_axis_tlast   (siAPP_Tcp_Data_tlast),
    .s_axis_tready  (siAPP_Tcp_Data_tready),
    //-- To NTS ------------------------
    .m_axis_tdata   (soNTS_Tcp_Data_tdata),
    .m_axis_tkeep   (soNTS_Tcp_Data_tkeep),
    .m_axis_tlast   (soNTS_Tcp_Data_tlast),
    .m_axis_tvalid  (soNTS_Tcp_Data_tvalid),
    .m_axis_tready  (soNTS_Tcp_Data_tready)
  );
  
  AxisRegisterSlice_16 APP_NTS_Tcp_Meta (
    .aclk           (piClk),
    .aresetn        (~piRst),
    //-- From APP ----------------------
    .s_axis_tdata   (siAPP_Tcp_Meta_tdata),
    .s_axis_tvalid  (siAPP_Tcp_Meta_tvalid),
    .s_axis_tready  (siAPP_Tcp_Meta_tready),
    //-- To NTS ------------------------
    .m_axis_tdata   (soNTS_Tcp_Meta_tdata),
    .m_axis_tvalid  (soNTS_Tcp_Meta_tvalid),
    .m_axis_tready  (soNTS_Tcp_Meta_tready)
  );
   
  AxisRegisterSlice_24 NTS_APP_Tcp_DSts (
    .aclk           (piClk),
    .aresetn        (~piRst),
    //-- From NTS ----------------------
    .s_axis_tdata   (siNTS_Tcp_DSts_tdata),
    .s_axis_tvalid  (siNTS_Tcp_DSts_tvalid),
    .s_axis_tready  (siNTS_Tcp_DSts_tready),
    //-- To APP ------------------------
    .m_axis_tdata   (soAPP_Tcp_DSts_tdata),
    .m_axis_tvalid  (soAPP_Tcp_DSts_tvalid),
    .m_axis_tready  (soAPP_Tcp_DSts_tready)
  );
    
  //------------------------------------------------------
  //-- TAIF / Rx Data Interfaces 
  //------------------------------------------------------
  AxisRegisterSlice_64 NTS_APP_Tcp_Data (
    .aclk           (piClk),
    .aresetn        (~piRst),
    //-- From NTS ----------------------
    .s_axis_tdata   (siNTS_Tcp_Data_tdata),
    .s_axis_tvalid  (siNTS_Tcp_Data_tvalid),
    .s_axis_tkeep   (siNTS_Tcp_Data_tkeep),
    .s_axis_tlast   (siNTS_Tcp_Data_tlast),
    .s_axis_tready  (siNTS_Tcp_Data_tready),
    //-- To APP ------------------------
    .m_axis_tdata   (soAPP_Tcp_Data_tdata),
    .m_axis_tkeep   (soAPP_Tcp_Data_tkeep),
    .m_axis_tlast   (soAPP_Tcp_Data_tlast),
    .m_axis_tvalid  (soAPP_Tcp_Data_tvalid),
    .m_axis_tready  (soAPP_Tcp_Data_tready)
  );
        
  AxisRegisterSlice_16 NTS_APP_Tcp_Meta (
    .aclk           (piClk),
    .aresetn        (~piRst),
    //-- From NTS ----------------------
    .s_axis_tdata   (siNTS_Tcp_Meta_tdata),
    .s_axis_tvalid  (siNTS_Tcp_Meta_tvalid),
    .s_axis_tready  (siNTS_Tcp_Meta_tready),
    //-- To APP ------------------------
    .m_axis_tdata   (soAPP_Tcp_Meta_tdata),
    .m_axis_tvalid  (soAPP_Tcp_Meta_tvalid),
    .m_axis_tready  (soAPP_Tcp_Meta_tready)
  );

  AxisRegisterSlice_104 NTS_APP_Tcp_Notif (
    .aclk           (piClk),
    .aresetn        (~piRst),
    //-- From NTS ----------------------
    .s_axis_tdata   (siNTS_Tcp_Notif_tdata),
    .s_axis_tvalid  (siNTS_Tcp_Notif_tvalid),
    .s_axis_tready  (siNTS_Tcp_Notif_tready),
    //-- To APP ------------------------
    .m_axis_tdata   (soAPP_Tcp_Notif_tdata),
    .m_axis_tvalid  (soAPP_Tcp_Notif_tvalid),
    .m_axis_tready  (soAPP_Tcp_Notif_tready)
  );
  
  AxisRegisterSlice_32 APP_NTS_Tcp_DReq (
    .aclk           (piClk),
    .aresetn        (~piRst),
    //-- From APP ----------------------
    .s_axis_tdata   (siAPP_Tcp_DReq_tdata),
    .s_axis_tvalid  (siAPP_Tcp_DReq_tvalid),
    .s_axis_tready  (siAPP_Tcp_DReq_tready),
    //-- To NTS ------------------------
    .m_axis_tdata   (soNTS_Tcp_DReq_tdata),
    .m_axis_tvalid  (soNTS_Tcp_DReq_tvalid),
    .m_axis_tready  (soNTS_Tcp_DReq_tready)
  );
  
  //------------------------------------------------------
  //-- TAIF / Tx Ctlr Interfaces
  //------------------------------------------------------
  AxisRegisterSlice_48 APP_NTS_Tcp_OpnReq (
    .aclk           (piClk),
    .aresetn        (~piRst),
    //-- From APP ----------------------
    .s_axis_tdata   (siAPP_Tcp_OpnReq_tdata),
    .s_axis_tvalid  (siAPP_Tcp_OpnReq_tvalid),
    .s_axis_tready  (siAPP_Tcp_OpnReq_tready),
    //-- To NTS ------------------------
    .m_axis_tdata   (soNTS_Tcp_OpnReq_tdata),
    .m_axis_tvalid (soNTS_Tcp_OpnReq_tvalid),
    .m_axis_tready  (soNTS_Tcp_OpnReq_tready)
  );  
  
  AxisRegisterSlice_24 NTS_APP_Tcp_OpnRep (
   .aclk           (piClk),
   .aresetn        (~piRst),
   //-- From NTS ----------------------
   .s_axis_tdata   (siNTS_Tcp_OpnRep_tdata),
   .s_axis_tvalid  (siNTS_Tcp_OpnRep_tvalid),
   .s_axis_tready  (siNTS_Tcp_OpnRep_tready),
   //-- To APP ------------------------
   .m_axis_tdata   (soAPP_Tcp_OpnRep_tdata),
   .m_axis_tvalid (soAPP_Tcp_OpnRep_tvalid),
   .m_axis_tready  (soAPP_Tcp_OpnRep_tready)
 );
 
 AxisRegisterSlice_16 APP_NTS_Tcp_ClsReq (
   .aclk           (piClk),
   .aresetn        (~piRst),
   //-- From APP ----------------------
   .s_axis_tdata   (siAPP_Tcp_ClsReq_tdata),
   .s_axis_tvalid  (siAPP_Tcp_ClsReq_tvalid),
   .s_axis_tready  (siAPP_Tcp_ClsReq_tready),
   //-- To NTS ------------------------
   .m_axis_tdata   (soNTS_Tcp_ClsReq_tdata),
   .m_axis_tvalid (soNTS_Tcp_ClsReq_tvalid),
   .m_axis_tready  (soNTS_Tcp_ClsReq_tready)
 );
  
  //------------------------------------------------------
  //-- TAIF / Rx Ctlr Interfaces 
  //------------------------------------------------------
  AxisRegisterSlice_16 APP_NTS_Tcp_LsnReq (
   .aclk           (piClk),
   .aresetn        (~piRst),
   //-- From APP ----------------------
   .s_axis_tdata   (siAPP_Tcp_LsnReq_tdata),
   .s_axis_tvalid  (siAPP_Tcp_LsnReq_tvalid),
   .s_axis_tready  (siAPP_Tcp_LsnReq_tready),
   //-- To NTS ------------------------
   .m_axis_tdata   (soNTS_Tcp_LsnReq_tdata),
   .m_axis_tvalid (soNTS_Tcp_LsnReq_tvalid),
   .m_axis_tready  (soNTS_Tcp_LsnReq_tready)
 );
  
 AxisRegisterSlice_8 NTS_APP_Tcp_LsnRep (
  .aclk           (piClk),
  .aresetn        (~piRst),
  //-- From NTS ----------------------
  .s_axis_tdata   (siNTS_Tcp_LsnRep_tdata),
  .s_axis_tvalid  (siNTS_Tcp_LsnRep_tvalid),
  .s_axis_tready  (siNTS_Tcp_LsnRep_tready),
  //-- To APP ------------------------
  .m_axis_tdata   (soAPP_Tcp_LsnRep_tdata),
  .m_axis_tvalid  (soAPP_Tcp_LsnRep_tvalid),
  .m_axis_tready  (soAPP_Tcp_LsnRep_tready)
); 

endmodule
