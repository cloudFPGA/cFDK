/*******************************************************************************
 * Copyright 2016 -- 2021 IBM Corporation
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *******************************************************************************/

// *****************************************************************************
// *
// *                             cloudFPGA
// *
// *----------------------------------------------------------------------------
// *
// * Title : Flash version of the the 10G Ethernet I/F instantiated by the SHELL. 
// *
// * File    : tenGigEth_Flash.v
// *
// * Created : Dec. 2017
// * Authors : Francois Abel <fab@zurich.ibm.com>
// *
// * Devices : xcku060-ffva1156-2-i
// * Tools   : Vivado v2016.4 (64-bit)
// * Depends : None
// *
// * Description : This is the toplevel design for the 10 Gigabit Ethernet I/F
// *    instantiated by the shell of the FMKU2595 module equipped with a XCKU60
// *    device. It is referred to as the Flash version because it integrates a  
// *    loopback turn between the network layers L2 and L3 of the ETH0 interface.
// *    When this loopback is enabled, the data output by the AXI4-S interface
// *    of ETH0 are passed back to the AXI4-S input of the same ETH0. Otherwise,
// *    this module is neutral and data pass through it untouched.  
// * 
// * Parameters:
// *
// * Comments:
// *
// *****************************************************************************


// *****************************************************************************
// **  ETH0 - 10G ETHERNET WITH LOOPBACK TURN
// *****************************************************************************

module TenGigEth_Flash (

  //-- Clocks and Resets inputs ------------------
  input             piTOP_156_25Clk,    // Freerunning
  input             piCLKT_Gt_RefClk_n,
  input             piCLKT_Gt_RefClk_p,
  input             piTOP_Reset,

  //-- Clocks and Resets outputs -----------------
  output            poSHL_CoreClk,
  output            poSHL_CoreResetDone,

   //-- MMIO : Control inputs and Status outputs -
  input             piMMIO_RxEqualizerMode,
  input  [ 3:0]     piMMIO_TxDriverSwing,
  input  [ 4:0]     piMMIO_TxPreCursor,
  input  [ 4:0]     piMMIO_TxPostCursor,
  input             piMMIO_PcsLoopbackEn,
  input             piMMIO_MacLoopbackEn,
  input             piMMIO_MacAddrSwapEn,
  output            poMMIO_CoreReady,
  output            poMMIO_QpllLock,

  //-- ECON : Gigabit Transceivers ---------------
  input             piECON_Gt_n,
  input             piECON_Gt_p,
  output            poECON_Gt_n,
  output            poECON_Gt_p,
   
  //-- NTS : Network-Transport-Session -----------
  //---- Input AXI-Write Stream Interface --------
  input     [63:0]  siLY3_Data_tdata,
  input     [7:0]   siLY3_Data_tkeep,
  input             siLY3_Data_tlast,
  input             siLY3_Data_tvalid,
  output            siLY3_Data_tready,
  //-- LY3 : Output Axi-Wirte Stream Interface ---
  output     [63:0] soLY3_Data_tdata,
  output     [7:0]  soLY3_Data_tkeep,
  output            soLY3_Data_tlast,
  output            soLY3_Data_tvalid,
   input            soLY3_Data_tready
  
); // End of PortList
   
// *****************************************************************************


  //============================================================================
  //  SIGNAL DECLARATIONS
  //============================================================================

  //-- Clocks and Resets --------------------------
  wire        sETH_CoreResetDone;
  wire        sETH_CoreClk;  // Generated by the ETHernet core. 
                             // Use it to clock the TX datapath.

  //-- AXI4 Stream ETH0 < -> NTS0 -----------------
  wire [63:0] ssETH_ELP_Data_tdata,  ssELP_ETH_Data_tdata;
  wire [ 7:0] ssETH_ELP_Data_tkeep,  ssELP_ETH_Data_tkeep;
  wire        ssETH_ELP_Data_tvalid, ssELP_ETH_Data_tvalid;
  wire        ssETH_ELP_Data_tlast,  ssELP_ETH_Data_tlast;
  wire        ssETH_ELP_Data_tready, ssELP_ETH_Data_tready;
    
  //-- End of signal declarations ---------------


  //============================================================================
  //  INST ETH: 10G ETHERNET SUBSYSTEM (OSI Network Layers 1+2)
  //============================================================================
  TenGigEth ETH (
    
    //-- Clocks and Resets inputs ----------------
    .piTOP_156_25Clk              (piTOP_156_25Clk),    // Freerunning
    .piCLKT_Gt_RefClk_n           (piCLKT_Gt_RefClk_n),
    .piCLKT_Gt_RefClk_p           (piCLKT_Gt_RefClk_p),
    .piTOP_Reset                  (piTOP_Reset),
      
    //-- Clocks and Resets outputs ---------------
    .poSHL_CoreClk                (sETH_CoreClk),
    .poSHL_CoreResetDone          (sETH_CoreResetDone),
       
    //-- MMIO : Control inputs and Status outputs 
    .piMMIO_RxEqualizerMode       (piMMIO_RxEqualizerMode),
    .piMMIO_TxDriverSwing         (piMMIO_TxDriverSwing),
    .piMMIO_TxPreCursor           (piMMIO_TxPreCursor),
    .piMMIO_TxPostCursor          (piMMIO_TxPostCursor),
    .piMMIO_PcsLoopbackEn         (piMMIO_PcsLoopbackEn),
    .poMMIO_CoreReady             (poMMIO_CoreReady),
    .poMMIO_QpllLock              (poMMIO_QpllLock),
    
    //-- ECON : Gigabit Transceivers -------------
    .piECON_Gt_n                  (piECON_Gt_n),
    .piECON_Gt_p                  (piECON_Gt_p),
    .poECON_Gt_n                  (poECON_Gt_n),
    .poECON_Gt_p                  (poECON_Gt_p),
         
    //-- LY3 : Layer-3 Input Interface -----------
    .siLY3_Data_tdata             (ssELP_ETH_Data_tdata),
    .siLY3_Data_tkeep             (ssELP_ETH_Data_tkeep),
    .siLY3_Data_tlast             (ssELP_ETH_Data_tlast),
    .siLY3_Data_tvalid            (ssELP_ETH_Data_tvalid),
    .siLY3_Data_tready            (ssELP_ETH_Data_tready),
 
    //-- LY3 : Layer-3 Output Interface ----------
    .soLY3_Data_tdata             (ssETH_ELP_Data_tdata),
    .soLY3_Data_tkeep             (ssETH_ELP_Data_tkeep),
    .soLY3_Data_tlast             (ssETH_ELP_Data_tlast),
    .soLY3_Data_tvalid            (ssETH_ELP_Data_tvalid),
    .soLY3_Data_tready            (ssETH_ELP_Data_tready)
  
  );  // End of PortList
    

  //============================================================================
  //  INST ELP: ETHERNET LOOPBACK TURN
  //============================================================================
  TenGigEth_Loop ELP (
      
    //-- Clocks and Resets inputs ----------------
    .piETH_CoreClk          (sETH_CoreClk),
    .piETH_CoreResetDone    (sETH_CoreResetDone),
    
    // -- MMIO : Ctrl Inp and Status Out ---------
    .piMMIO_LoopbackEn      (piMMIO_MacLoopbackEn),
    .piMMIO_AddrSwapEn      (piMMIO_MacAddrSwapEn),

     //-- LY2 : Input AXI-Write Stream Interface -
    .siLY2_Data_tdata       (ssETH_ELP_Data_tdata),
    .siLY2_Data_tkeep       (ssETH_ELP_Data_tkeep),
    .siLY2_Data_tlast       (ssETH_ELP_Data_tlast),
    .siLY2_Data_tvalid      (ssETH_ELP_Data_tvalid),
    .siLY2_Data_tready      (ssETH_ELP_Data_tready),
    
    // LY2 : Input AXI-Write Stream Interface ----
    .soLY2_Data_tdata       (ssELP_ETH_Data_tdata),
    .soLY2_Data_tkeep       (ssELP_ETH_Data_tkeep),
    .soLY2_Data_tlast       (ssELP_ETH_Data_tlast),
    .soLY2_Data_tvalid      (ssELP_ETH_Data_tvalid),
    .soLY2_Data_tready      (ssELP_ETH_Data_tready),
    
    //-- LY3 : Input AXI-Write Stream Interface --
    .siLY3_Data_tdata       (siLY3_Data_tdata),
    .siLY3_Data_tkeep       (siLY3_Data_tkeep),
    .siLY3_Data_tlast       (siLY3_Data_tlast),
    .siLY3_Data_tvalid      (siLY3_Data_tvalid),
    .siLY3_Data_tready      (siLY3_Data_tready),
    
    // LY3 : Input AXI-Write Stream Interface ----
    .soLY3_Data_tdata       (soLY3_Data_tdata),
    .soLY3_Data_tkeep       (soLY3_Data_tkeep),
    .soLY3_Data_tlast       (soLY3_Data_tlast),
    .soLY3_Data_tvalid      (soLY3_Data_tvalid),
    .soLY3_Data_tready      (soLY3_Data_tready)
                  
  );


  //============================================================================
  //  COMB: CONTINUOUS OUTPUT PORT ASSIGNMENTS
  //============================================================================
  assign poSHL_CoreClk       = sETH_CoreClk;
  assign poSHL_CoreResetDone = sETH_CoreResetDone;

endmodule
