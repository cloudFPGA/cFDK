//                              -*- Mode: Verilog -*-
// *****************************************************************************
// *
// *                             cloudFPGA
// *            All rights reserved -- Property of IBM
// *
// *----------------------------------------------------------------------------
// *
// * Title : UDP Application Register Slice (UARS)
// *
// * Created : Apr. 2020
// * Authors : Francois Abel <fab@zurich.ibm.com>
// *
// * Tools   : Vivado v2016.4 (64-bit)
// * Depends : None
// *
// * Description : A placeholder containing the Axis Register Slice (ARS) 
// *    components involved in the UDP application interface of the Network
// *    Transport Stack (NTS). The use of such an Axis register slice is not
// *    a prerequisit but it is used here to provide timing isolation and to
// *    ease the place and routing phase.
// *
// *          +-----+     +----+     +---+
// *          |     <-----+    <-----+   |
// *          | NTS |     |UARS|     |APP|
// *          |     +----->    +----->   |
// *          +-----+     +----+     +---+
// *
// *****************************************************************************

`timescale 1ns / 1ps

// *****************************************************************************
// **  MODULE - UDP APPLICATION REGISTER SLICE
// *****************************************************************************

module UdpApplicationRegisterSlice

(

  //------------------------------------------------------
  //-- This is typically the Global Clock used all over the SHELL
  //------------------------------------------------------ 
  input           piClk,
  
  //------------------------------------------------------
  //-- This is typically the Global Reset used by the entire SHELL
  //--  or the OSI-Layer-5 reset generated by the MMIO. 
  //------------------------------------------------------ 
  input           piRst,
 
  //------------------------------------------------------
  //-- APP / Udp / Tx Data Interfaces (.i.e APP->UARS)
  //------------------------------------------------------
  //---- Axis4-Stream UDP Data ---------------
  input  [ 63:0]  siAPP_Udp_Data_tdata ,
  input  [  7:0]  siAPP_Udp_Data_tkeep ,
  input           siAPP_Udp_Data_tlast ,
  input           siAPP_Udp_Data_tvalid,
  output          siAPP_Udp_Data_tready,
  //---- Axis4-Stream UDP Metadata -----------
  input   [95:0]  siAPP_Udp_Meta_tdata ,
  input           siAPP_Udp_Meta_tvalid,
  output          siAPP_Udp_Meta_tready,
  //---- Axis4Stream UDP Data Length ---------
  input   [15:0]  siAPP_Udp_DLen_tdata ,
  input           siAPP_Udp_DLen_tvalid,
  output          siAPP_Udp_DLen_tready,
    
  //------------------------------------------------------
  //-- APP / Udp / Rx Data Interfaces (.i.e UARS-->APP)
  //------------------------------------------------------
  //---- Axis4-Stream UDP Data ---------------
  output  [63:0]  soAPP_Udp_Data_tdata ,
  output  [ 7:0]  soAPP_Udp_Data_tkeep ,
  output          soAPP_Udp_Data_tlast ,
  output          soAPP_Udp_Data_tvalid,
  input           soAPP_Udp_Data_tready,
  //---- Axis4-Stream UDP Metadata -----------
  output  [95:0]  soAPP_Udp_Meta_tdata ,
  output          soAPP_Udp_Meta_tvalid,
  input           soAPP_Udp_Meta_tready,
  
  //------------------------------------------------------
  //-- APP / Udp / Rx Ctrl Interfaces (.i.e UARS<-->APP)
  //------------------------------------------------------
  //---- Axis4-Stream UDP Listen Request -----
  input   [15:0]  siAPP_Udp_LsnReq_tdata ,
  input           siAPP_Udp_LsnReq_tvalid,
  output          siAPP_Udp_LsnReq_tready,
  //---- Axis4-Stream UDP Listen Reply --------
  output  [ 7:0]  soAPP_Udp_LsnRep_tdata ,
  output          soAPP_Udp_LsnRep_tvalid,
  input           soAPP_Udp_LsnRep_tready,
  //---- Axis4-Stream UDP Close Request ------
  input   [15:0]  siAPP_Udp_ClsReq_tdata ,
  input           siAPP_Udp_ClsReq_tvalid,
  output          siAPP_Udp_ClsReq_tready,
  //---- Axis4-Stream UDP Close Reply ---------
  output  [ 7:0]  soAPP_Udp_ClsRep_tdata ,
  output          soAPP_Udp_ClsRep_tvalid,
  input           soAPP_Udp_ClsRep_tready,

  //------------------------------------------------------
  //-- NTS / Udp / Tx Data Interfaces (.i.e UARS-->NTS)
  //------------------------------------------------------
  //---- Axis4-Stream UDP Data ---------------
  output [ 63:0]  soNTS_Udp_Data_tdata ,
  output [  7:0]  soNTS_Udp_Data_tkeep ,
  output          soNTS_Udp_Data_tlast ,
  output          soNTS_Udp_Data_tvalid,
  input           soNTS_Udp_Data_tready,
  //---- Axis4-Stream UDP Metadata -----------
  output  [95:0]  soNTS_Udp_Meta_tdata ,
  output          soNTS_Udp_Meta_tvalid,
  input           soNTS_Udp_Meta_tready,
  //---- Axis4Stream UDP Data Length ---------
  output  [15:0]  soNTS_Udp_DLen_tdata ,
  output          soNTS_Udp_DLen_tvalid,
  input           soNTS_Udp_DLen_tready,
    
  //------------------------------------------------------
  //-- NTS / Udp / Rx Data Interfaces (.i.e NTS<-->UARS)
  //------------------------------------------------------
  //---- Axis4-Stream UDP Data ---------------
  input   [63:0]  siNTS_Udp_Data_tdata ,
  input   [ 7:0]  siNTS_Udp_Data_tkeep ,
  input           siNTS_Udp_Data_tlast ,
  input           siNTS_Udp_Data_tvalid,
  output          siNTS_Udp_Data_tready,
  //---- Axis4-Stream UDP Metadata -----------
  input   [95:0]  siNTS_Udp_Meta_tdata ,
  input           siNTS_Udp_Meta_tvalid,
  output          siNTS_Udp_Meta_tready,
  
  //------------------------------------------------------
  //-- NTS / Udp / Rx Ctrl Interfaces (.i.e NTS<-->UARS)
  //------------------------------------------------------
  //---- Axis4-Stream UDP Listen Request -----
  output  [15:0]  soNTS_Udp_LsnReq_tdata ,
  output          soNTS_Udp_LsnReq_tvalid,
  input           soNTS_Udp_LsnReq_tready,
  //---- Axis4-Stream UDP Listen Reply --------
  input   [ 7:0]  siNTS_Udp_LsnRep_tdata ,
  input           siNTS_Udp_LsnRep_tvalid,
  output          siNTS_Udp_LsnRep_tready,
  //---- Axis4-Stream UDP Close Request ------
  output  [15:0]  soNTS_Udp_ClsReq_tdata ,
  output          soNTS_Udp_ClsReq_tvalid,
  input           soNTS_Udp_ClsReq_tready,
  //---- Axis4-Stream UDP Listen Reply --------
  input   [ 7:0]  siNTS_Udp_ClsRep_tdata ,
  input           siNTS_Udp_ClsRep_tvalid,
  output          siNTS_Udp_ClsRep_tready
  
);  // End of PortList


  // *****************************************************************************
  // **  STRUCTURE
  // *****************************************************************************
   
  //------------------------------------------------------
  //-- UAIF / Tx Data Interfaces
  //------------------------------------------------------ 
  AxisRegisterSlice_64 APP_NTS_Udp_Data (
    .aclk           (piClk),
    .aresetn        (~piRst),
    //-- From APP ----------------------
    .s_axis_tdata  (siAPP_Udp_Data_tdata) ,
    .s_axis_tkeep  (siAPP_Udp_Data_tkeep) ,
    .s_axis_tlast  (siAPP_Udp_Data_tlast) ,
    .s_axis_tvalid (siAPP_Udp_Data_tvalid),
    .s_axis_tready (siAPP_Udp_Data_tready),     
    //-- To NTS ------------------------
    .m_axis_tdata  (soNTS_Udp_Data_tdata) ,
    .m_axis_tkeep  (soNTS_Udp_Data_tkeep) ,
    .m_axis_tlast  (soNTS_Udp_Data_tlast) ,
    .m_axis_tvalid (soNTS_Udp_Data_tvalid),
    .m_axis_tready (soNTS_Udp_Data_tready)
  );

  AxisRegisterSlice_96 APP_NTS_Udp_Meta (
    .aclk           (piClk),
    .aresetn        (~piRst),
    //-- From NTS ----------------------
    .s_axis_tdata  (siAPP_Udp_Meta_tdata) ,
    .s_axis_tvalid (siAPP_Udp_Meta_tvalid),
    .s_axis_tready (siAPP_Udp_Meta_tready),     
    //-- To APP ------------------------
    .m_axis_tdata  (soNTS_Udp_Meta_tdata) ,
    .m_axis_tvalid (soNTS_Udp_Meta_tvalid),
    .m_axis_tready (soNTS_Udp_Meta_tready)
  );  
   
  AxisRegisterSlice_16 APP_NTS_Udp_DLen (
    .aclk           (piClk),
    .aresetn        (~piRst),
    //-- From NTS ----------------------
    .s_axis_tdata  (siAPP_Udp_DLen_tdata) ,
    .s_axis_tvalid (siAPP_Udp_DLen_tvalid),
    .s_axis_tready (siAPP_Udp_DLen_tready),     
    //-- To APP ------------------------
    .m_axis_tdata  (soNTS_Udp_DLen_tdata) ,
    .m_axis_tvalid (soNTS_Udp_DLen_tvalid),
    .m_axis_tready (soNTS_Udp_DLen_tready)
  );
    
  //------------------------------------------------------
  //-- UAIF / Rx Data Interfaces
  //------------------------------------------------------
  AxisRegisterSlice_64 NTS_APP_Udp_Data (
    .aclk           (piClk),
    .aresetn        (~piRst),
    //-- From NTS ----------------------
    .s_axis_tdata  (siNTS_Udp_Data_tdata) ,
    .s_axis_tkeep  (siNTS_Udp_Data_tkeep) ,
    .s_axis_tlast  (siNTS_Udp_Data_tlast) ,
    .s_axis_tvalid (siNTS_Udp_Data_tvalid),
    .s_axis_tready (siNTS_Udp_Data_tready),     
    //-- To APP ------------------------
    .m_axis_tdata  (soAPP_Udp_Data_tdata) ,
    .m_axis_tkeep  (soAPP_Udp_Data_tkeep) ,
    .m_axis_tlast  (soAPP_Udp_Data_tlast) ,
    .m_axis_tvalid (soAPP_Udp_Data_tvalid),
    .m_axis_tready (soAPP_Udp_Data_tready)
  );
  
  AxisRegisterSlice_96 NTS_APP_Udp_Meta (
    .aclk           (piClk),
    .aresetn        (~piRst),
    //-- From NTS ----------------------
    .s_axis_tdata  (siNTS_Udp_Meta_tdata) ,
    .s_axis_tvalid (siNTS_Udp_Meta_tvalid),
    .s_axis_tready (siNTS_Udp_Meta_tready),     
    //-- To APP ------------------------
    .m_axis_tdata  (soAPP_Udp_Meta_tdata) ,
    .m_axis_tvalid (soAPP_Udp_Meta_tvalid),
    .m_axis_tready (soAPP_Udp_Meta_tready)
  );
  
  //------------------------------------------------------
  //-- UAIF / Rx Ctrl Interfaces (.i.e NTS-->APP)
  //------------------------------------------------------  
  AxisRegisterSlice_16 NTS_APP_Udp_LsnReq (
    .aclk           (piClk),
    .aresetn        (~piRst),
    //-- From NTS ----------------------
    .s_axis_tdata  (siAPP_Udp_LsnReq_tdata) ,
    .s_axis_tvalid (siAPP_Udp_LsnReq_tvalid),
    .s_axis_tready (siAPP_Udp_LsnReq_tready),     
    //-- To APP ------------------------
    .m_axis_tdata  (soNTS_Udp_LsnReq_tdata) ,
    .m_axis_tvalid (soNTS_Udp_LsnReq_tvalid),
    .m_axis_tready (soNTS_Udp_LsnReq_tready)
  );

  AxisRegisterSlice_8 NTS_APP_Udp_LsnRep (
    .aclk           (piClk),
    .aresetn        (~piRst),
    //-- From NTS ----------------------
    .s_axis_tdata  (siNTS_Udp_LsnRep_tdata) ,
    .s_axis_tvalid (siNTS_Udp_LsnRep_tvalid),
    .s_axis_tready (siNTS_Udp_LsnRep_tready),     
    //-- To APP ------------------------
    .m_axis_tdata  (soAPP_Udp_LsnRep_tdata) ,
    .m_axis_tvalid (soAPP_Udp_LsnRep_tvalid),
    .m_axis_tready (soAPP_Udp_LsnRep_tready)
  );
  
  AxisRegisterSlice_16 NTS_APP_Udp_ClsReq (
    .aclk           (piClk),
    .aresetn        (~piRst),
    //-- From NTS ----------------------
    .s_axis_tdata  (siAPP_Udp_ClsReq_tdata) ,
    .s_axis_tvalid (siAPP_Udp_ClsReq_tvalid),
    .s_axis_tready (siAPP_Udp_ClsReq_tready),     
    //-- To APP ------------------------
    .m_axis_tdata  (soNTS_Udp_ClsReq_tdata) ,
    .m_axis_tvalid (soNTS_Udp_ClsReq_tvalid),
    .m_axis_tready (soNTS_Udp_ClsReq_tready)
  );
  
  AxisRegisterSlice_8 NTS_APP_Udp_ClsRep (
      .aclk           (piClk),
      .aresetn        (~piRst),
      //-- From NTS ----------------------
      .s_axis_tdata  (siNTS_Udp_ClsRep_tdata) ,
      .s_axis_tvalid (siNTS_Udp_ClsRep_tvalid),
      .s_axis_tready (siNTS_Udp_ClsRep_tready),     
      //-- To APP ------------------------
      .m_axis_tdata  (soAPP_Udp_ClsRep_tdata) ,
      .m_axis_tvalid (soAPP_Udp_ClsRep_tvalid),
      .m_axis_tready (soAPP_Udp_ClsRep_tready)
    );

endmodule
