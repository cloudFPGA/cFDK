// *****************************************************************************
// *
// *                             cloudFPGA
// *            All rights reserved -- Property of IBM
// *
// *----------------------------------------------------------------------------
// *
// * Title : Flash version of the the 10G Ethernet I/F instantiated by the SHELL. 
// *
// * File    : tenGigEth_Flash.v
// *
// * Created : Dec. 2017
// * Authors : Francois Abel <fab@zurich.ibm.com>
// *
// * Devices : xcku060-ffva1156-2-i
// * Tools   : Vivado v2016.4 (64-bit)
// * Depends : None
// *
// * Description : This is the toplevel design for the 10 Gigabit Ethernet I/F
// *    instantiated by the shell of the FMKU2595 module equipped with a XCKU60
// *    device. It is referred to as the Flash version because it integrates a  
// *    loopback turn between the network layers L2 and L3 of the ETH0 interface.
// *    When this loopback is enabled, the data output by the AXI4-S interface
// *    of ETH0 are passed back to the AXI4-S input of the same ETH0. Otherwise,
// *    this module is neutral and data pass through it untouched.  
// * 
// * Parameters:
// *
// * Comments:
// *
// *****************************************************************************


// *****************************************************************************
// **  ETH0 - 10G ETHERNET WITH LOOPBACK TURN
// *****************************************************************************

module TenGigEth_Flash (

  //-- Clocks and Resets inputs ------------------
  input             piTOP_156_25Clk,    // Freerunning
  input             piCLKT_Gt_RefClk_n,
  input             piCLKT_Gt_RefClk_p,
  input             piTOP_Reset,

  //-- Clocks and Resets outputs -----------------
  output            poETH0_CoreClk,
  output            poETH0_CoreResetDone,

  //-- MMIO : Ctrl inputs and Status outputs -----
  input             piMMIO_Eth0_RxEqualizerMode,
  input             piMMIO_Eth0_PcsLoopbackEn,
  input             piMMIO_Eth0_MacLoopbackEn,
  input             piMMIO_Eth0_MacAddrSwapEn,
  output            poETH0_Mmio_CoreReady,
  output            poETH0_Mmio_QpllLock,
  output            poETH0_Mmio_ResetDone,

  //-- ECON : Gigabit Transceivers ---------------
  input             piECON_Eth0_Gt_n,
  input             piECON_Eth0_Gt_p,
  output            poETH0_Econ_Gt_n,
  output            poETH0_Econ_Gt_p,
   
  //-- LY3 : Input AXI-Write Stream Interface ----
  input     [63:0]  piLY3_Eth0_Axis_tdata,
  input     [7:0]   piLY3_Eth0_Axis_tkeep,
  input             piLY3_Eth0_Axis_tlast,
  input             piLY3_Eth0_Axis_tvalid,
  output            poETH0_Ly3_Axis_tready,
  
  //-- LY3 : Output Axi-Wirte Stream Interface ---
  input             piLY3_Eth0_Axis_tready,
  output     [63:0] poETH0_Ly3_Axis_tdata,
  output     [7:0]  poETH0_Ly3_Axis_tkeep,
  output            poETH0_Ly3_Axis_tlast,
  output            poETH0_Ly3_Axis_tvalid
  
); // End of PortList
   
// *****************************************************************************


  //============================================================================
  //  SIGNAL DECLARATIONS
  //============================================================================

  //-- Clocks and Resets --------------------------
  wire        sETH0_CoreResetDone;
  wire        sETH0_CoreClk;  // Generated by the ETH core. 
                              // Use it to clock the TX datapath.

  //-- AXI4 Stream ETH0 < -> NTS0 -----------------
  wire [63:0] sETH_Elp_Axis_tdata,  sELP_Eth_Axis_tdata;
  wire [ 7:0] sETH_Elp_Axis_tkeep,  sELP_Eth_Axis_tkeep;
  wire        sETH_Elp_Axis_tvalid, sELP_Eth_Axis_tvalid;
  wire        sETH_Elp_Axis_tlast,  sELP_Eth_Axis_tlast;
  wire        sELP_Eth_Axis_tready, sETH_Elp_Axis_tready;
    
  //-- End of signal declarations ---------------


  //============================================================================
  //  INST ETH: 10G ETHERNET SUBSYSTEM (OSI Network Layers 1+2)
  //============================================================================
  TenGigEth ETH (
    
    //-- Clocks and Resets inputs ----------------
    .piTOP_156_25Clk              (piTOP_156_25Clk),    // Freerunning
    .piCLKT_Gt_RefClk_n           (piCLKT_Gt_RefClk_n),
    .piCLKT_Gt_RefClk_p           (piCLKT_Gt_RefClk_p),
    .piTOP_Reset                  (piTOP_Reset),
      
    //-- Clocks and Resets outputs ---------------
    .poETH0_CoreClk               (sETH0_CoreClk),
    .poETH0_CoreResetDone         (sETH0_CoreResetDone),
       
    //-- MMIO : Control inputs and Status outputs 
    .piMMIO_Eth0_RxEqualizerMode  (piMMIO_Eth0_RxEqualizerMode),
    .piMMIO_Eth0_PcsLoopbackEn    (piMMIO_Eth0_PcsLoopbackEn),
    .poETH0_Mmio_CoreReady        (poETH0_Mmio_CoreReady),
    .poETH0_Mmio_QpllLock         (poETH0_Mmio_QpllLock),
    
    //-- ECON : Gigabit Transceivers -------------
    .piECON_Eth0_Gt_n             (piECON_Eth0_Gt_n),
    .piECON_Eth0_Gt_p             (piECON_Eth0_Gt_p),
    .poETH0_Econ_Gt_n             (poETH0_Econ_Gt_n),
    .poETH0_Econ_Gt_p             (poETH0_Econ_Gt_p),
         
    //-- LY3 : Input AXI-Write Stream Interface --
    .piLY3_Eth0_Axis_tdata        (sELP_Eth_Axis_tdata),
    .piLY3_Eth0_Axis_tkeep        (sELP_Eth_Axis_tkeep),
    .piLY3_Eth0_Axis_tlast        (sELP_Eth_Axis_tlast),
    .piLY3_Eth0_Axis_tvalid       (sELP_Eth_Axis_tvalid),
    .poETH0_Ly3_Axis_tready       (sETH_Elp_Axis_tready),

    //-- LY3 : Output AXI-Write Stream Interface -
    .piLY3_Eth0_Axis_tready       (sELP_Eth_Axis_tready),
    .poETH0_Ly3_Axis_tdata        (sETH_Elp_Axis_tdata),
    .poETH0_Ly3_Axis_tkeep        (sETH_Elp_Axis_tkeep),
    .poETH0_Ly3_Axis_tlast        (sETH_Elp_Axis_tlast),
    .poETH0_Ly3_Axis_tvalid       (sETH_Elp_Axis_tvalid)
  
  );
    

  //============================================================================
  //  INST ELP: ETHERNET LOOPBACK TURN
  //============================================================================
  TenGigEth_Loop ELP (
      
        //-- Clocks and Resets inputs ------------
        .piETH0_CoreClk         (sETH0_CoreClk),
        .piETH0_CoreResetDone   (sETH0_CoreResetDone),
      
        // -- MMIO : Ctrl Inp and Status Out -----
        .piMMIO_LoopbackEn      (piMMIO_Eth0_MacLoopbackEn),
        .piMMIO_AddrSwapEn      (piMMIO_Eth0_MacAddrSwapEn),

         //-- LY2 : Input AXI-Write Stream Interface ----
        .piLY2_Elp_Axis_tdata   (sETH_Elp_Axis_tdata),
        .piLY2_Elp_Axis_tkeep   (sETH_Elp_Axis_tkeep),
        .piLY2_Elp_Axis_tlast   (sETH_Elp_Axis_tlast),
        .piLY2_Elp_Axis_tvalid  (sETH_Elp_Axis_tvalid),
        .poELP_Ly2_Axis_tready  (sELP_Eth_Axis_tready),
        
        // LY2 : Input AXI-Write Stream Interface ------
        .piLY2_Elp_Axis_tready  (sETH_Elp_Axis_tready),
        .poELP_Ly2_Axis_tdata   (sELP_Eth_Axis_tdata),
        .poELP_Ly2_Axis_tkeep   (sELP_Eth_Axis_tkeep),
        .poELP_Ly2_Axis_tlast   (sELP_Eth_Axis_tlast),
        .poELP_Ly2_Axis_tvalid  (sELP_Eth_Axis_tvalid),
        
        //-- LY3 : Input AXI-Write Stream Interface ----
        .piLY3_Elp_Axis_tdata   (piLY3_Eth0_Axis_tdata),
        .piLY3_Elp_Axis_tkeep   (piLY3_Eth0_Axis_tkeep),
        .piLY3_Elp_Axis_tlast   (piLY3_Eth0_Axis_tlast),
        .piLY3_Elp_Axis_tvalid  (piLY3_Eth0_Axis_tvalid),        
        .poELP_Ly3_Axis_tready  (poETH0_Ly3_Axis_tready),
        
        // LY3 : Input AXI-Write Stream Interface ------
        .piLY3_Elp_Axis_tready  (piLY3_Eth0_Axis_tready),
        .poELP_Ly3_Axis_tdata   (poETH0_Ly3_Axis_tdata),
        .poELP_Ly3_Axis_tkeep   (poETH0_Ly3_Axis_tkeep),
        .poELP_Ly3_Axis_tlast   (poETH0_Ly3_Axis_tlast),
        .poELP_Ly3_Axis_tvalid  (poETH0_Ly3_Axis_tvalid)
                      
      );


  //============================================================================
  //  COMB: CONTINUOUS OUTPUT PORT ASSIGNMENTS
  //============================================================================
  assign poETH0_CoreClk       = sETH0_CoreClk;
  assign poETH0_CoreResetDone = sETH0_CoreResetDone;

endmodule
